class Register;
    string name;
    rand bit [3:0] name;