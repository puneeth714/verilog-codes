//and_gate using gate_level modeling
module and_gate(a,b,c);
//a,b are inputs and c is output
input a;
input b;
output c;
 and(c,a,b);
endmodule
//end and gate

