module andd(
    a,b,c,d
);
    
endmodule