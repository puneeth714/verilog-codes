module tb;
string ex="Good morning";
intial begin
$display("%s",ex);
end
endmodule
