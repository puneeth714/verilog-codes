module four_bit_full_adder(a[0:3],b[0:3],c[0:3],d[0:4]);
input a[0:3],b[0:3],c[0:3];
output d[0:4];
endmodule
