module full_adder(a,b,c);
input a;
input b;
output c;
endmodule
