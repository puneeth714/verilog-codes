module while_loop()